library IEEE;
use IEEE.std_logic_1164.all;

entity ALU_Total is 
  port (
    A : in std_logic_vector(31 downto 0);
    B : in std_logic_vector(31 downto 0);
    ALU_Control : in std_logic_vector(3 downto 0);
    Branch_Control : in std_logic_vector(2 downto 0);
    S : out std_logic_vector(31 downto 0);
    zero : out std_logic;
    overflow : out std_logic
  );
end ALU_Total;

architecture structural of ALU_Total is 
  -- 0000 AND, 0001 OR, 0011 XOR
  -- 0010 ADD, 0110 SUB 
  -- 0100 SLL, 0101 SRL, 0111 SRA, 1000 SLT
  -- 1011 LUI

  signal s_AND, s_OR, s_XOR : std_logic_vector(31 downto 0);
  signal s_AddSub : std_logic_vector(31 downto 0);
  signal s_controlAdder : std_logic;
  signal s_C, s_Overflw : std_logic;
  signal s_BarrelShifted : std_logic_vector(31 downto 0);
  signal s_zero : std_logic;
  signal s_setLessThan : std_logic_vector(31 downto 0);

  component AddSub_overflow is 
    generic(N : integer := 16);
    port (
      A_i : in  std_logic_vector(N-1 downto 0);
      B_i : in  std_logic_vector(N-1 downto 0);
      nAdd_Sub : in  std_logic;  -- 0 => Add, 1 => Subtract
      S_i : out std_logic_vector(N-1 downto 0);
      C_out : out std_logic;
      Overflow_out : out std_logic
    );
  end component;

  component mux_16t1 is 
    generic (WIDTH : integer := 32);
    port (
        sel    : in  std_logic_vector(3 downto 0);
        in0    : in  std_logic_vector(WIDTH-1 downto 0);
        in1    : in  std_logic_vector(WIDTH-1 downto 0);
        in2    : in  std_logic_vector(WIDTH-1 downto 0);
        in3    : in  std_logic_vector(WIDTH-1 downto 0);
        in4    : in  std_logic_vector(WIDTH-1 downto 0);
        in5    : in  std_logic_vector(WIDTH-1 downto 0);
        in6    : in  std_logic_vector(WIDTH-1 downto 0);
        in7    : in  std_logic_vector(WIDTH-1 downto 0);
        in8    : in  std_logic_vector(WIDTH-1 downto 0);
        in9    : in  std_logic_vector(WIDTH-1 downto 0);
        in10   : in  std_logic_vector(WIDTH-1 downto 0);
        in11   : in  std_logic_vector(WIDTH-1 downto 0);
        in12   : in  std_logic_vector(WIDTH-1 downto 0);
        in13   : in  std_logic_vector(WIDTH-1 downto 0);
        in14   : in  std_logic_vector(WIDTH-1 downto 0);
        in15   : in  std_logic_vector(WIDTH-1 downto 0);
        y      : out std_logic_vector(WIDTH-1 downto 0)
    );
  end component;

  component barrel_shifter is 
   port (
    data_in     : in  std_logic_vector(31 downto 0);
    shift_amt    : in  std_logic_vector(4 downto 0);
    ALU_Control : in std_logic_vector(3 downto 0);
    result    : out std_logic_vector(31 downto 0)
  );
  end component;

  component Branch is
    port (
      Difference : in std_logic_vector(31 downto 0);
      Branch_Control : in std_logic_vector(2 downto 0);
      C_out : in std_logic;
      Overflow : in std_logic;
      Zero : out std_logic
    );
  end component;

begin 
  s_AND <= A and B;
  s_OR <= A or B;
  s_XOR <= A xor B;

  s_controlAdder <= '1' when (ALU_Control = "0110" or 
				ALU_Control = "1000" or 
				ALU_Control = "1001" ) else '0';

  adder : AddSub_overflow 
    generic map (N => 32)
    port map (
      A_i => A,
      B_i => B,
      nAdd_Sub => s_controlAdder,
      S_i => s_AddSub,
      C_out => s_C,
      Overflow_out => s_Overflw 
    );
    
  shifty_time : barrel_shifter 
    port map (
      data_in => A,
      shift_amt => B(4 downto 0),
      ALU_Control => ALU_Control,
      result => s_BarrelShifted
    );

  branch_time : Branch 
    port map (
      Difference => s_AddSub,
      Branch_Control => Branch_Control,
	C_out => s_C,
      Overflow => s_Overflw,
      Zero => s_zero
    );

zero <= s_zero;

s_setLessThan <= x"00000001" when (s_zero = '1') else x"00000000";

  big_mux : mux_16t1
    generic map (WIDTH => 32)
    port map (
      sel => ALU_Control,
      in0 => s_AND,
      in1 => s_OR,
      in2 => s_AddSub,
      in3 => s_XOR,
      in4 => s_BarrelShifted,
      in5 => s_BarrelShifted,
      in6 => s_AddSub,
      in7 => s_BarrelShifted,
      in8 => s_setLessThan,
      in9 => s_setLessThan,
      in10 => s_BarrelShifted,
      in11 => B,
      in12 => x"00000000",
      in13 => x"00000000",
      in14 => x"00000000",
      in15 => x"00000000",
      y => S
    );

    overflow <= '1' when (s_Overflw = '1' and (ALU_Control = "0010" or ALU_Control = "0110")) else '0';
    

end structural;
