-- Zevan Gustafson
-- zevang@iastate.edu

-- mux2t1.vhd with structural iplementation

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity mux2t1 is 
port(i_D0 : in std_logic;
	i_D1 : in std_logic;
	i_S : in std_logic;
	o_O : out std_logic);
end mux2t1;

-- Structural
architecture behavior of mux2t1 is

signal wire1, wire2, wire3 : std_logic;

component andg2 is
port(i_A : in std_logic;
	i_B : in std_logic;
	o_F : out std_logic);
end component;

component org2 is 
port (i_A : in std_logic;
	i_B : in std_logic;
	o_F : out std_logic);
end component;

component invg is 
port (i_A : in std_logic;
	o_F : out std_logic);
end component;

begin

not_gate1 : invg 
port map ( i_A => i_S,
	o_F => wire1);

and_gate1 : andg2
port map ( i_A => wire1,
	i_B => i_D0,
	o_F => wire2);

and_gate2 : andg2
port map ( i_A => i_S,
	i_B => i_D1,
	o_F => wire3);

or_gate1 : org2
port map ( i_A => wire2,
	i_B => wire3,
	o_F => o_O);

end behavior;
