-- Test bench for mux2t1_N
-- Zevan Gustafson zevang@iastate.edu

