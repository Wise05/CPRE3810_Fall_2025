library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity tb_ALU_Total is
  generic(gCLK_HPER   : time := 50 ns;
          N : integer := 32);
end tb_ALU_Total;

architecture behavior of tb_ALU_Total is
  
  -- Calculate the clock period as twice the half-period
  constant cCLK_PER  : time := gCLK_HPER * 2;


  component ALU_Total
     port ( 
    	A : in std_logic_vector(31 downto 0);
     	B : in std_logic_vector(31 downto 0);
     	ALU_Control : in std_logic_vector(3 downto 0);
     	Branch_Control : in std_logic_vector(2 downto 0);
     	S : out std_logic_vector(31 downto 0);
     	zero : out std_logic;
     	overflow : out std_logic
);
  end component;

signal s_CLK : std_logic := '0';  
signal s_A : std_logic_vector(31 downto 0) := (others => '0');
  signal s_B : std_logic_vector(31 downto 0) := (others => '0');
  signal s_ALU_Control : std_logic_vector(3 downto 0) := (others => '0');
  signal s_Branch_Control : std_logic_vector(2 downto 0) := (others => '0');
  signal s_S : std_logic_vector(31 downto 0) := (others => '0');
  signal s_zero : std_logic := '0';
  signal s_overflow : std_logic := '0';

begin

  DUT: ALU_Total
  port map(
    	   A => s_A,
    	   B => s_B,
    	   ALU_Control => s_ALU_Control,
   	   Branch_Control => s_Branch_Control,
    	   S => s_S,
    	   zero => s_zero,
    	   overflow => s_overflow
);
	

  P_CLK: process
  begin
    s_CLK <= '0';
    wait for gCLK_HPER;
    s_CLK <= '1';
    wait for gCLK_HPER;
  end process;

  P_TB: process
  begin

-- add, sub, and, or, xor, sll, sra, beq, bne, blt

--1 Add
    s_A <= "00000000000000000000000000000000";
    s_B <= "00000000000000000000000000000001";
    s_ALU_Control <= "0010";
    s_Branch_Control <= "000";
    wait for cCLK_PER; 

--2 Sub
    s_A <= "00000000000000000000000000000001";
    s_B <= "00000000000000000000000000000001";
    s_ALU_Control <= "0110";
    s_Branch_Control <= "000";
    wait for cCLK_PER; 

--3 And
    s_A <= "00000000000000000000000000000001";
    s_B <= "00000000000000000000000000000000";
    s_ALU_Control <= "0000";
    s_Branch_Control <= "000";
    wait for cCLK_PER; 

--4 Or
    s_A <= "00000000000000000000000000000001";
    s_B <= "00000000000000000000000000000000";
    s_ALU_Control <= "0001";
    s_Branch_Control <= "000";
    wait for cCLK_PER; 

--5 Xor
    s_A <= "00000000000000000000000000000001";
    s_B <= "00000000000000000000000000000001";
    s_ALU_Control <= "0011";
    s_Branch_Control <= "000";
    wait for cCLK_PER; 

--6 Sll
    s_A <= "00000000000000000000000000000001";
    s_B <= "00000000000000000000000000000001";
    s_ALU_Control <= "0100";
    s_Branch_Control <= "000";
    wait for cCLK_PER; 

--7 Sra
    s_A <= "00000000000000000000000000000001";
    s_B <= "00000000000000000000000000000001";
    s_ALU_Control <= "0111";
    s_Branch_Control <= "000";
    wait for cCLK_PER; 

--8 Beq
    s_A <= "00000000000000000000000000000001";
    s_B <= "00000000000000000000000000000001";
    s_ALU_Control <= "0110";
    s_Branch_Control <= "000";
    wait for cCLK_PER; 

--9 Bne
    s_A <= "00000000000000000000000000000001";
    s_B <= "00000000000000000000000000000000";
    s_ALU_Control <= "0110";
    s_Branch_Control <= "001";
    wait for cCLK_PER; 

--10 Blt
    s_A <= "00000000000000000000000000000010";
    s_B <= "00000000000000000000000000000001";
    s_ALU_Control <= "0110";
    s_Branch_Control <= "010";
    wait for cCLK_PER; 

    wait;
  end process;
  
end behavior;
