-- Zevan Gustafson
-- dffg_N
-- N bit register file

library IEEE;
use IEEE.std_logic_1161.all;

entity dffg_N is 
    generic(N : integer := 32);
    port(i_CLK        : in std_logic;
       i_RST        : in std_logic;     -- Reset input
       i_WE         : in std_logic;     -- Write enable input
       i_D          : in std_logic_vector(N-1 downto 0);     -- Data value input
       o_Q          : out std_logic_vector(N-1 downto 0)); -- Data value output
end dffg_N;

architecture structural of dffg_N is

    component dffg is 
        port(i_CLK        : in std_logic;     -- Clock input
        i_RST        : in std_logic;     -- Reset input
        i_WE         : in std_logic;     -- Write enable input
        i_D          : in std_logic;     -- Data value input
        o_Q          : out std_logic);
    end component;

begin

    G_NBIT_REGISTER: for i in 0 to N-1 generate
        REGI: dffg port map (
            i_CLK => i_CLK,
            iRST => iRST,
            i_WE => iWE,
            iD => iD(i),
            o_Q => o_Q(i)
        );
    end generate G_NBIT_REGISTER;

end structural;


