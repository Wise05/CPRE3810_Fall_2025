library IEEE;
use IEEE.std_logic_1164.all;


entity MEM_WB is --13 inputs
  port (
    in_dmem         : in std_logic_vector(31 downto 0);
    in_MemtoReg     : in std_logic;
    in_RegWrite     : in std_logic;
    in_regWrite_addr : in std_logic_vector(4 downto 0);
    in_mux          : in std_logic_vector(31 downto 0);
    in_alu          : in std_logic_vector(31 downto 0);
    in_load         : in std_logic_vector(2 downto 0);
    in_halt         : in std_logic;
    WE              : in std_logic;
    out_dmem        : out std_logic_vector(31 downto 0);
    out_MemtoReg    : out std_logic;
    out_RegWrite    : out std_logic;
    out_regWrite_addr : out std_logic_vector(4 downto 0);
    out_mux         : out std_logic_vector(31 downto 0);
    out_alu         : out std_logic_vector(31 downto 0);
    out_load        : out std_logic_vector(2 downto 0);
    out_halt        : out std_logic;
    RST             : in std_logic;
    CLK             : in std_logic
  );
end MEM_WB;


architecture structural of MEM_WB is 
  
  component Nbit_reg is 
    generic(N : integer := 32); 
    port (
        in_1 : in std_logic_vector(N-1 downto 0);
	WE : in std_logic;
	out_1 : out std_logic_vector(N-1 downto 0);
	RST : in std_logic;
	CLK: in std_logic
);
  end component;

begin

dmem_reg: Nbit_reg
	generic map (N => 32)
	port map (
		in_1 => in_dmem,
		WE => WE,
		out_1 => out_dmem,
		RST => RST,
		CLK => CLK
    );

MemtoReg_reg: Nbit_reg
	generic map (N => 1)
	port map (
		in_1(0) => in_MemtoReg,
		WE => WE,
		out_1(0) => out_MemtoReg,
		RST => RST,
		CLK => CLK
    );
    
RegWrite_reg: Nbit_reg
	generic map (N => 1)
	port map (
		in_1(0) => in_RegWrite,
		WE => WE,
		out_1(0) => out_RegWrite,
		RST => RST,
		CLK => CLK
    );

RegWriteAddress_reg: Nbit_reg
  generic map (N => 5)
  port map (
	in_1 => in_regWrite_addr,
	WE => WE,
	out_1 => out_regWrite_addr,
	RST => RST,
	CLK => CLK
    );

load_reg : Nbit_reg
  generic map (N => 3)
  port map (
	in_1 => in_load,
	WE => WE,
	out_1 => out_load,
	RST => RST,
	CLK => CLK
    );

halt_reg: Nbit_reg
	generic map (N => 1)
	port map (
		in_1(0) => in_halt,
		WE => WE,
		out_1(0) => out_halt,
		RST => RST,
		CLK => CLK
    );
    
mux_reg: Nbit_reg
	generic map (N => 32)
	port map (
		in_1 => in_mux,
		WE => WE,
		out_1 => out_mux,
		RST => RST,
		CLK => CLK
    );

alu_reg: Nbit_reg
	generic map (N => 32)
	port map (
		in_1 => in_alu,
		WE => WE,
		out_1 => out_alu,
		RST => RST,
		CLK => CLK
    );

end structural;
