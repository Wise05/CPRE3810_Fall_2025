-- tb N-bit one's complementor
-- Zephaniah Gustafson

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_textio.all;  -- For logic types I/O
library std;
use std.textio.all;

entity tb_ones_comp_N is
generic (gCLK_HPER : time := 10 ns;
	DATA_WIDTH : integer := 32);
end tb_ones_comp_N;

architecture mixed of tb_ones_comp_N is 

component ones_comp_N is 
generic (N : integer := 32);
port(i_C : in std_logic_vector(N-1 downto 0);
	o_C : out std_logic_vector(N-1 downto 0));
end component;

signal si_C : std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
signal so_C : std_logic_vector(DATA_WIDTH-1 downto 0);

begin 

DUT0: ones_comp_N
generic map (N => DATA_WIDTH)
port map(
	i_C => si_C,
	o_C => so_C);

P_TEST_CASES: process
begin 
wait for gCLK_HPER/2;

-- Test case 1:
si_C <= x"00000000";
wait for gCLK_HPER * 2;
-- expect so_C = FFFFFFFF

-- Test case 2:
si_C <= x"12341234";
wait for gCLK_HPER * 2;
-- expect so_C = EDCBEDCB

-- Test case 3:
si_C <= x"CAFEF00D";
wait for gCLK_HPER * 2;
-- expect so_C = 35010FF2;

wait;
end process;
end mixed;
-- 