-- library IEEE;
-- use IEEE.stad_logic_1164.all;
-- 
 entity ALU_Total is 
--   port (
--     A : in std_logic_vector(31 downto 0);
--     B : in std_logic_vector(31 downto 0);
--     ALU_Control : in std_logic_vector(3 downto 0);
--     Branch_Control : in std_logic_vector(2 downto 0);
--     S : out std_logic_vector(31 downto 0);
--     zero : out std_logic;
--     overflow : out std_logic;
--   );
 end ALU_Total;
 
 architecture structural of ALU_Total is 
--   -- 0000 AND, 0001 OR, 0011 XOR
--   -- 0010 ADD, 0110 SUB 
--   -- 0100 SLL, 0101 SRL, 0111 SRA, 1000 SLT
-- 
--   signal s_AND, s_OR, s_XOR : std_logic_vector(31 downto 0);
--   signal s_AddSub : std_logic_vector(31 downto 0);
--   signal s_BarrelShifted : std_logic_vector(31 downto 0);
-- 
--   component add_sub_N is 
--     generic(N : integer := 16);
--     port (
--       A_i : in  std_logic_vector(N-1 downto 0);
--       B_i : in  std_logic_vector(N-1 downto 0);
--       nAdd_Sub : in  std_logic;  -- 0 => Add, 1 => Subtract
--       S_i : out std_logic_vector(N-1 downto 0);
--       C_out : out std_logic
--     );
--   end component;
-- 
--   component mux_16t1 is 
--     generic (WIDTH : integer := 32);
--     port (
--         sel    : in  std_logic_vector(3 downto 0);
--         in0    : in  std_logic_vector(WIDTH-1 downto 0);
--         in1    : in  std_logic_vector(WIDTH-1 downto 0);
--         in2    : in  std_logic_vector(WIDTH-1 downto 0);
--         in3    : in  std_logic_vector(WIDTH-1 downto 0);
--         in4    : in  std_logic_vector(WIDTH-1 downto 0);
--         in5    : in  std_logic_vector(WIDTH-1 downto 0);
--         in6    : in  std_logic_vector(WIDTH-1 downto 0);
--         in7    : in  std_logic_vector(WIDTH-1 downto 0);
--         in8    : in  std_logic_vector(WIDTH-1 downto 0);
--         in9    : in  std_logic_vector(WIDTH-1 downto 0);
--         in10   : in  std_logic_vector(WIDTH-1 downto 0);
--         in11   : in  std_logic_vector(WIDTH-1 downto 0);
--         in12   : in  std_logic_vector(WIDTH-1 downto 0);
--         in13   : in  std_logic_vector(WIDTH-1 downto 0);
--         in14   : in  std_logic_vector(WIDTH-1 downto 0);
--         in15   : in  std_logic_vector(WIDTH-1 downto 0);
--         y      : out std_logic_vector(WIDTH-1 downto 0)
--     );
--   end component;
-- 
--   component BarrelShifter is 
--     
--   end component;
-- 
--   component BranchController is
--     PC : in std_logic_vector(31 downto 0);
--     offset : in std_logic_vector(31 downto 0);
--     difference : in std_logic_vector(31 downto 0);
--   end component;
 begin 
--   s_AND <= A and B;
--   s_OR <= A or B;
--   s_XOR <= A xor B;
-- 
-- 
end structural;
