library IEEE;
use IEEE.std_logic_1164.all;
use work.regfile_pkg.all;

entity fetch is 
  -- inputs jump, branch, immediate (extended), zero flag
  port (
      
 )
