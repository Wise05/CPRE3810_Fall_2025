library IEEE;
use IEEE.std_logic_1164.all;

entity dffg is
  port(
    i_CLK : in std_logic;
    i_RST : in std_logic;
    i_WE  : in std_logic;
    i_D   : in std_logic;
    o_Q   : out std_logic
  );
end entity;

architecture behavioral of dffg is
  signal r_Q : std_logic := '0';  
begin
  process(i_CLK, i_RST)
  begin
    if i_RST = '1' then
      r_Q <= '0'; 
    elsif rising_edge(i_CLK) then
      if i_WE = '1' then
        r_Q <= i_D;
      end if;
    end if;
  end process;

  o_Q <= r_Q;
end architecture;

