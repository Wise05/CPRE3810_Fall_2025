-- Zevan Gustafson zevang@iastate.edu

-- mux2t1_dataflow test bench
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_textio.all;  -- For logic types I/O
library std;
--use std.env.all;                -- For hierarchical/external signals
use std.textio.all; 

entity tb_mux2t1_dataflow is 
	generic (gCLK_HPER : time := 10 ns);
end tb_mux2t1_dataflow;

architecture mixed of tb_mux2t1_dataflow is 

constant cCLK_PER : time := gCLK_HPER * 2;

component mux2t1_dataflow is 
	port (i_D0 : in std_logic;
	i_D1 : in std_logic;
	i_S : in std_logic;
	o_O : out std_logic);
end component;

signal CLK : std_logic := '0';
signal D0 : std_logic := '0';
signal D1 : std_logic := '0';
signal S : std_logic := '0';
signal O : std_logic;

begin

DUT0: mux2t1_dataflow
port map(
	i_D0 => D0,
	i_D1 => D1,
	i_S => S,
	o_O => O);

P_CLK: process
  begin
    CLK <= '1';         -- clock starts at 1
    wait for gCLK_HPER; -- after half a cycle
    CLK <= '0';         -- clock becomes a 0 (negative edge)
    wait for gCLK_HPER; -- after half a cycle, process begins evaluation again
  end process; 

P_TEST_CASES: process
  begin
    wait for gCLK_HPER/2; -- for waveform clarity, I prefer not to change inputs on clk edges

    -- Test case 1:
D0 <= '0';
D1 <= '0';
S <= '0';
wait for gCLK_HPER*2;

    -- Test case 2:
D0 <= '0';
D1 <= '0';
S <= '1';
wait for gCLK_HPER*2;

-- Test case 3
D0 <= '0';
D1 <= '1';
S <= '0';
wait for gCLK_HPER*2;

-- Test case 4 
D0 <= '0';
D1 <= '1';
S <= '1';
wait for gCLK_HPER*2;

-- Test case 5
D0 <= '1';
D1 <= '0';
S <= '0';
wait for gCLK_HPER*2;

-- Test case 6
D0 <= '1';
D1 <= '0';
S <= '1';
wait for gCLK_HPER*2;

-- Test case 7
D0 <= '1';
D1 <= '1';
S <= '0';
wait for gCLK_HPER*2;

-- Test case 8
D0 <= '1';
D1 <= '1';
S <= '1';
wait for gCLK_HPER*2;

    wait;
  end process;

end mixed;